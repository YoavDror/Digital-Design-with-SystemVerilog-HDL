`timescale 1ns/1ps

module hello_world;
  initial begin
    $display("Hello World!");
  end
endmodule
